2803:6780::/32
167.249.20.0/22
132.255.208.0/22
